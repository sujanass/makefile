//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////Copyright © 2022 Vivartan Technologies., All rights reserved////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                              //
//All works published under Zilla_Gen_0 by Vivartan Technologies is copyrighted by the Association and ownership// 
//of all right, title and interest in and to the works remains with Vivartan Technologies. No works or documents//
//published under Zilla_Gen_0 by Vivartan Technologies may be reproduced,transmitted or copied without the expre//
//-ss written permission of Vivartan Technologies will be considered as a violations of Copyright Act and it may//
//lead to legal action.                                                                                         //
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/*////////////////////////////////////////////////////////////////////////////////////////////////////////////////
* File Name : riscv_package.svh

* Purpose : package for riscv

* Creation Date : 17-03-2023

* Last Modified : Thu 04 May 2023 01:13:17 PM IST

* Created By :  sharon
*/

package test_package;
    import uvm_pkg::*;

    `include "uvm_macros.svh"

    //test
    `include "./../test/riscv_base_test.svh"
    `include "./../test/riscv_inst_test.svh"
    `include "./../test/riscv_sb_inst_test.svh"
    `include "./../test/riscv_i_inst_test.svh"

  
  
  endpackage
    


